package types_pkg;

  typedef enum {ADD, SUB, MUL, DIV} op_type;

endpackage: types_pkg
